/*
    Copyright 2020 UCLouvain

    Licensed under the Solderpad Hardware Licence, Version 2.0 (the "License");
    you may not use this file except in compliance with the License.
    You may obtain a copy of the License at

        https://solderpad.org/licenses/SHL-2.0/

    Unless required by applicable law or agreed to in writing, software
    distributed under the License is distributed on an "AS IS" BASIS,
    WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
    See the License for the specific language governing permissions and
    limitations under the License.
*/

(* fv_prop = "_mux", fv_strat = "assumed", fv_order = d *)
module MSKmux #(parameter d=1) (sel, in_true, in_false, out);

	(* fv_type = "control" *) input sel;
	(* fv_type = "sharing", fv_latency = 0 *) input  [d-1:0] in_true;
	(* fv_type = "sharing", fv_latency = 0 *) input  [d-1:0] in_false;
	(* fv_type = "sharing", fv_latency = 0 *) output [d-1:0] out;

	assign out = sel ? in_true : in_false;

endmodule
