/*
    Copyright 2020 UCLouvain

    Licensed under the Solderpad Hardware Licence, Version 2.0 (the "License");
    you may not use this file except in compliance with the License.
    You may obtain a copy of the License at

        https://solderpad.org/licenses/SHL-2.0/

    Unless required by applicable law or agreed to in writing, software
    distributed under the License is distributed on an "AS IS" BASIS,
    WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
    See the License for the specific language governing permissions and
    limitations under the License.
*/
/*
    This module implements the xtime operation used to 
    generate the 32-bits constants.
*/
module xtime
(
    input [31:0] x_in,
    output [31:0] x_out
);

wire [31:0] b = (x_in >> 31);
assign x_out = (x_in << 1) ^ b ^(b << 8);

endmodule
