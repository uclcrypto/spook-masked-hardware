/*
    Copyright 2020 UCLouvain

    Licensed under the Solderpad Hardware Licence, Version 2.0 (the "License");
    you may not use this file except in compliance with the License.
    You may obtain a copy of the License at

        https://solderpad.org/licenses/SHL-2.0/

    Unless required by applicable law or agreed to in writing, software
    distributed under the License is distributed on an "AS IS" BASIS,
    WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
    See the License for the specific language governing permissions and
    limitations under the License.
*/
/*
    This module creates a valid sharing for non-sensitive value.
    It uses 0 instead of randomness to create the shares. 
*/
(* fv_prop = "affine", fv_strat = "assumed", fv_order = d *)
module cst_mask #(parameter d=1, parameter count=1) (cst, out);

	(* fv_type = "control" *)       input [count-1:0] cst;
	(* fv_type = "sharing", fv_count = count, fv_latency = 0 *) output [count*d-1:0] out;

	genvar i;
	for(i=0; i<count; i=i+1) begin: i_gen_m
		assign out[i*d +: d] = { cst[i], {(d-1){1'b0}}};
	end

endmodule
